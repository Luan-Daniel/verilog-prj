library verilog;
use verilog.vl_types.all;
entity mux2x1_tb is
end mux2x1_tb;
