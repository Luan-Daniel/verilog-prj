/**
 * lab4
 * Aluno: Luan Daniel de Oliveira Melo (20102096)
 *
 ** lab4\src\half_adder.v **
 * Define um modulo para um meio somador de N bits
 */

module half_adder
#(parameter N = 4)
(a, b, s, c);
	input [N-1:0] a, b;
	output [N-1:0] s;
	output c;

	assign {c, s} = a + b;

endmodule //half_adder
