library verilog;
use verilog.vl_types.all;
entity half_adder_tb is
end half_adder_tb;
